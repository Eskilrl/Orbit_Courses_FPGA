module AND(
    //place inputs and outputs here:

    //Example:

    //input a,
    //input b,

    //output c
);


//Write your logic here:

    
endmodule